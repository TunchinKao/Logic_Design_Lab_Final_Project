//
//
//
//

`define c1 32'd261
`define c1_u 32'd277
`define d1_d 32'd277
`define d1 32'd293 
`define d1_u 32'd311
`define e1_d 32'd311
`define e1 32'd329
`define f1 32'd349
`define f1_u 32'd370
`define g1_d 32'd370
`define g1 32'd392
`define g1_u 32'd415
`define a1_d 32'd415
`define a1 32'd440
`define a1_u 32'd466
`define b1_d 32'd466
`define b1 32'd494
`define non 32'd20000 //slience (over freq.)

module Music (
	input [11:0] ibeatNum,	
	input [3:0] state,
	input [1:0] pitch,
	output reg [31:0] tone
);

reg [31:0] toneH, toneM, toneL;

always @(*) begin
	case (ibeatNum)		// 1/4 beat
		12'd0: toneH = `a1<<1;
		12'd1: toneH = `g1_u << 1;
		12'd2: toneH = `g1<<1;
		12'd3: toneH = `f1_u << 1;
		12'd4: toneH = `a1<<1;
		12'd5: toneH = `f1<<1;
		12'd6: toneH = `g1_d << 1;
		12'd7: toneH = `f1<<1;
		12'd8: toneH = `a1<<1;
		12'd9: toneH = `e1<<1;
		12'd10: toneH = `f1<<1;
		12'd11: toneH = `e1<<1;
		12'd12: toneH = `a1<<1;
		12'd13: toneH = `d1_u << 1;
		12'd14: toneH = `e1<<1;
		12'd15: toneH = `d1_u << 1;
		12'd16: toneH = `a1<<1;
		12'd17: toneH = `d1<<1;
		12'd18: toneH = `e1_d << 1;
		12'd19: toneH = `d1<<1;
		12'd20: toneH = `a1<<1;
		12'd21: toneH = `c1_u << 1;
		12'd22: toneH = `d1<<1;
		12'd23: toneH = `c1_u << 1;
		12'd24: toneH = `a1<<1;
		12'd25: toneH = `c1<<1;
		12'd26: toneH = `c1_u << 1;
		12'd27: toneH = `c1<<1;
		12'd28: toneH = `a1<<1;
		12'd29: toneH = `b1;
		12'd30: toneH = `c1<<1;
		12'd31: toneH = `b1;
		12'd32: toneH = `b1<<1;
		12'd33: toneH = `b1<<1;
		12'd34: toneH = `non;
		12'd35: toneH = `non;
		12'd36: toneH = `non;
		12'd37: toneH = `non;
		12'd38: toneH = `non;
		12'd39: toneH = `non;
		12'd40: toneH = `non;
		12'd41: toneH = `non;
		12'd42: toneH = `non;
		12'd43: toneH = `non;
		12'd44: toneH = `non;
		12'd45: toneH = `non;
		12'd46: toneH = `non;
		12'd47: toneH = `non;
		12'd48: toneH = `non;
		12'd49: toneH = `non;
		12'd50: toneH = `non;
		12'd51: toneH = `non;
		12'd52: toneH = `non;
		12'd53: toneH = `non;
		12'd54: toneH = `non;
		12'd55: toneH = `non;
		12'd56: toneH = `non;
		12'd57: toneH = `non;
		12'd58: toneH = `non;
		12'd59: toneH = `non;
		12'd60: toneH = `non;
		12'd61: toneH = `non;
		12'd62: toneH = `non;
		12'd63: toneH = `non;
		12'd64: toneH = `b1<<1;
		12'd65: toneH = `b1<<1;
		12'd66: toneH = `non;
		12'd67: toneH = `non;
		12'd68: toneH = `non;
		12'd69: toneH = `non;
		12'd70: toneH = `non;
		12'd71: toneH = `non;
		12'd72: toneH = `non;
		12'd73: toneH = `non;
		12'd74: toneH = `non;
		12'd75: toneH = `non;
		12'd76: toneH = `non;
		12'd77: toneH = `non;
		12'd78: toneH = `non;
		12'd79: toneH = `non;
		12'd80: toneH = `non;
		12'd81: toneH = `non;
		12'd82: toneH = `non;
		12'd83: toneH = `non;
		12'd84: toneH = `non;
		12'd85: toneH = `non;
		12'd86: toneH = `non;
		12'd87: toneH = `non;
		12'd88: toneH = `non;
		12'd89: toneH = `non;
		12'd90: toneH = `non;
		12'd91: toneH = `non;
		12'd92: toneH = `a1<<1;
		12'd93: toneH = `a1<<1;
		12'd94: toneH = `e1<<1;
		12'd95: toneH = `e1<<1;
		12'd96: toneH = `b1;
		12'd97: toneH = `b1;
		12'd98: toneH = `non;
		12'd99: toneH = `non;
		12'd100: toneH = `non;
		12'd101: toneH = `non;
		12'd102: toneH = `c1_u << 1;
		12'd103: toneH = `c1_u << 1;
		12'd104: toneH = `non;
		12'd105: toneH = `non;
		12'd106: toneH = `non;
		12'd107: toneH = `non;
		12'd108: toneH = `d1<<1;
		12'd109: toneH = `d1<<1;
		12'd110: toneH = `non;
		12'd111: toneH = `non;
		12'd112: toneH = `b1;
		12'd113: toneH = `b1;
		12'd114: toneH = `d1_d << 1;
		12'd115: toneH = `d1_d << 1;
		12'd116: toneH = `non;
		12'd117: toneH = `non;
		12'd118: toneH = `d1<<1;
		12'd119: toneH = `d1<<1;
		12'd120: toneH = `non;
		12'd121: toneH = `non;
		12'd122: toneH = `non;
		12'd123: toneH = `non;
		12'd124: toneH = `a1<<1;
		12'd125: toneH = `a1<<1;
		12'd126: toneH = `b1_d << 1;
		12'd127: toneH = `b1_d << 1;
		12'd128: toneH = `b1<<1;
		12'd129: toneH = `b1<<1;
		12'd130: toneH = `non;
		12'd131: toneH = `non;
		12'd132: toneH = `non;
		12'd133: toneH = `non;
		12'd134: toneH = `c1_u << 2;
		12'd135: toneH = `c1_u << 2;
		12'd136: toneH = `non;
		12'd137: toneH = `non;
		12'd138: toneH = `non;
		12'd139: toneH = `non;
		12'd140: toneH = `d1 << 2;
		12'd141: toneH = `d1 << 2;
		12'd142: toneH = `non;
		12'd143: toneH = `non;
		12'd144: toneH = `b1<<1;
		12'd145: toneH = `b1<<1;
		12'd146: toneH = `c1_u << 2;
		12'd147: toneH = `c1_u << 2;
		12'd148: toneH = `non;
		12'd149: toneH = `non;
		12'd150: toneH = `d1 << 2;
		12'd151: toneH = `d1 << 2;
		12'd152: toneH = `non;
		12'd153: toneH = `non;
		12'd154: toneH = `non;
		12'd155: toneH = `non;
		12'd156: toneH = `a1<<1;
		12'd157: toneH = `a1<<1;
		12'd158: toneH = `non;
		12'd159: toneH = `non;
		12'd160: toneH = `b1;
		12'd161: toneH = `b1;
		12'd162: toneH = `b1;
		12'd163: toneH = `b1;
		12'd164: toneH = `b1;
		12'd165: toneH = `b1;
		12'd166: toneH = `f1_u;
		12'd167: toneH = `f1_u;
		12'd168: toneH = `f1_u;
		12'd169: toneH = `f1_u;
		12'd170: toneH = `f1_u;
		12'd171: toneH = `f1_u;
		12'd172: toneH = `f1_u;
		12'd173: toneH = `f1_u;
		12'd174: toneH = `f1_u;
		12'd175: toneH = `f1_u;
		12'd176: toneH = `f1_u;
		12'd177: toneH = `f1_u;
		12'd178: toneH = `f1_u;
		12'd179: toneH = `f1_u;
		12'd180: toneH = `b1;
		12'd181: toneH = `b1;
		12'd182: toneH = `b1;
		12'd183: toneH = `b1;
		12'd184: toneH = `f1_u;
		12'd185: toneH = `f1_u;
		12'd186: toneH = `f1_u;
		12'd187: toneH = `f1_u;
		12'd188: toneH = `b1;
		12'd189: toneH = `b1;
		12'd190: toneH = `b1;
		12'd191: toneH = `b1;
		12'd192: toneH = `c1<<1;
		12'd193: toneH = `c1<<1;
		12'd194: toneH = `c1<<1;
		12'd195: toneH = `c1<<1;
		12'd196: toneH = `c1<<1;
		12'd197: toneH = `c1<<1;
		12'd198: toneH = `c1<<1;
		12'd199: toneH = `c1<<1;
		12'd200: toneH = `c1<<1;
		12'd201: toneH = `c1<<1;
		12'd202: toneH = `c1<<1;
		12'd203: toneH = `c1<<1;
		12'd204: toneH = `c1<<1;
		12'd205: toneH = `c1<<1;
		12'd206: toneH = `c1<<1;
		12'd207: toneH = `c1<<1;
		12'd208: toneH = `c1<<1;
		12'd209: toneH = `c1<<1;
		12'd210: toneH = `c1<<1;
		12'd211: toneH = `c1<<1;
		12'd212: toneH = `c1<<1;
		12'd213: toneH = `c1<<1;
		12'd214: toneH = `c1<<1;
		12'd215: toneH = `c1<<1;
		12'd216: toneH = `c1<<1;
		12'd217: toneH = `c1<<1;
		12'd218: toneH = `c1<<1;
		12'd219: toneH = `c1<<1;
		12'd220: toneH = `c1<<1;
		12'd221: toneH = `c1<<1;
		12'd222: toneH = `c1<<1;
		12'd223: toneH = `c1<<1;
		12'd224: toneH = `b1;
		12'd225: toneH = `b1;
		12'd226: toneH = `b1;
		12'd227: toneH = `b1;
		12'd228: toneH = `b1;
		12'd229: toneH = `b1;
		12'd230: toneH = `f1_u;
		12'd231: toneH = `f1_u;
		12'd232: toneH = `f1_u;
		12'd233: toneH = `f1_u;
		12'd234: toneH = `f1_u;
		12'd235: toneH = `f1_u;
		12'd236: toneH = `f1_u;
		12'd237: toneH = `f1_u;
		12'd238: toneH = `f1_u;
		12'd239: toneH = `f1_u;
		12'd240: toneH = `f1_u;
		12'd241: toneH = `f1_u;
		12'd242: toneH = `f1_u;
		12'd243: toneH = `f1_u;
		12'd244: toneH = `b1;
		12'd245: toneH = `b1;
		12'd246: toneH = `b1;
		12'd247: toneH = `b1;
		12'd248: toneH = `f1_u;
		12'd249: toneH = `f1_u;
		12'd250: toneH = `f1_u;
		12'd251: toneH = `f1_u;
		12'd252: toneH = `b1;
		12'd253: toneH = `b1;
		12'd254: toneH = `b1;
		12'd255: toneH = `b1;
		12'd256: toneH = `c1<<1;
		12'd257: toneH = `c1<<1;
		12'd258: toneH = `c1<<1;
		12'd259: toneH = `c1<<1;
		12'd260: toneH = `c1<<1;
		12'd261: toneH = `c1<<1;
		12'd262: toneH = `c1<<1;
		12'd263: toneH = `c1<<1;
		12'd264: toneH = `c1<<1;
		12'd265: toneH = `c1<<1;
		12'd266: toneH = `c1<<1;
		12'd267: toneH = `c1<<1;
		12'd268: toneH = `c1<<1;
		12'd269: toneH = `c1<<1;
		12'd270: toneH = `c1<<1;
		12'd271: toneH = `c1<<1;
		12'd272: toneH = `c1<<1;
		12'd273: toneH = `c1<<1;
		12'd274: toneH = `c1<<1;
		12'd275: toneH = `c1<<1;
		12'd276: toneH = `c1<<1;
		12'd277: toneH = `c1<<1;
		12'd278: toneH = `c1<<1;
		12'd279: toneH = `c1<<1;
		12'd280: toneH = `c1<<1;
		12'd281: toneH = `c1<<1;
		12'd282: toneH = `c1<<1;
		12'd283: toneH = `c1<<1;
		12'd284: toneH = `c1<<1;
		12'd285: toneH = `c1<<1;
		12'd286: toneH = `c1<<1;
		12'd287: toneH = `c1<<1;
		12'd288: toneH = `g1;
		12'd289: toneH = `g1;
		12'd290: toneH = `g1;
		12'd291: toneH = `g1;
		12'd292: toneH = `g1;
		12'd293: toneH = `g1;
		12'd294: toneH = `g1;
		12'd295: toneH = `g1;
		12'd296: toneH = `g1;
		12'd297: toneH = `g1;
		12'd298: toneH = `g1;
		12'd299: toneH = `g1;
		12'd300: toneH = `g1;
		12'd301: toneH = `g1;
		12'd302: toneH = `g1;
		12'd303: toneH = `g1;
		12'd304: toneH = `d1<<1;
		12'd305: toneH = `d1<<1;
		12'd306: toneH = `d1<<1;
		12'd307: toneH = `d1<<1;
		12'd308: toneH = `d1<<1;
		12'd309: toneH = `d1<<1;
		12'd310: toneH = `d1<<1;
		12'd311: toneH = `d1<<1;
		12'd312: toneH = `g1;
		12'd313: toneH = `g1;
		12'd314: toneH = `g1;
		12'd315: toneH = `g1;
		12'd316: toneH = `g1;
		12'd317: toneH = `g1;
		12'd318: toneH = `g1;
		12'd319: toneH = `g1;
		12'd320: toneH = `a1;
		12'd321: toneH = `a1;
		12'd322: toneH = `a1;
		12'd323: toneH = `a1;
		12'd324: toneH = `a1;
		12'd325: toneH = `a1;
		12'd326: toneH = `a1;
		12'd327: toneH = `a1;
		12'd328: toneH = `a1;
		12'd329: toneH = `a1;
		12'd330: toneH = `a1;
		12'd331: toneH = `a1;
		12'd332: toneH = `a1;
		12'd333: toneH = `a1;
		12'd334: toneH = `a1;
		12'd335: toneH = `a1;
		12'd336: toneH = `a1;
		12'd337: toneH = `a1;
		12'd338: toneH = `a1;
		12'd339: toneH = `a1;
		12'd340: toneH = `a1;
		12'd341: toneH = `a1;
		12'd342: toneH = `a1;
		12'd343: toneH = `a1;
		12'd344: toneH = `a1;
		12'd345: toneH = `a1;
		12'd346: toneH = `a1;
		12'd347: toneH = `a1;
		12'd348: toneH = `a1;
		12'd349: toneH = `a1;
		12'd350: toneH = `a1;
		12'd351: toneH = `a1;
		12'd352: toneH = `g1;
		12'd353: toneH = `g1;
		12'd354: toneH = `g1;
		12'd355: toneH = `g1;
		12'd356: toneH = `g1;
		12'd357: toneH = `g1;
		12'd358: toneH = `g1;
		12'd359: toneH = `g1;
		12'd360: toneH = `g1;
		12'd361: toneH = `g1;
		12'd362: toneH = `g1;
		12'd363: toneH = `g1;
		12'd364: toneH = `g1;
		12'd365: toneH = `g1;
		12'd366: toneH = `g1;
		12'd367: toneH = `g1;
		12'd368: toneH = `e1<<1;
		12'd369: toneH = `e1<<1;
		12'd370: toneH = `e1<<1;
		12'd371: toneH = `e1<<1;
		12'd372: toneH = `e1<<1;
		12'd373: toneH = `e1<<1;
		12'd374: toneH = `e1<<1;
		12'd375: toneH = `e1<<1;
		12'd376: toneH = `f1_u << 1;
		12'd377: toneH = `f1_u << 1;
		12'd378: toneH = `f1_u << 1;
		12'd379: toneH = `f1_u << 1;
		12'd380: toneH = `f1_u << 1;
		12'd381: toneH = `f1_u << 1;
		12'd382: toneH = `f1_u << 1;
		12'd383: toneH = `f1_u << 1;
		12'd384: toneH = `e1<<1;
		12'd385: toneH = `e1<<1;
		12'd386: toneH = `e1<<1;
		12'd387: toneH = `e1<<1;
		12'd388: toneH = `e1<<1;
		12'd389: toneH = `e1<<1;
		12'd390: toneH = `e1<<1;
		12'd391: toneH = `e1<<1;
		12'd392: toneH = `e1<<1;
		12'd393: toneH = `e1<<1;
		12'd394: toneH = `e1<<1;
		12'd395: toneH = `e1<<1;
		12'd396: toneH = `e1<<1;
		12'd397: toneH = `e1<<1;
		12'd398: toneH = `e1<<1;
		12'd399: toneH = `e1<<1;
		12'd400: toneH = `g1<<1;
		12'd401: toneH = `g1<<1;
		12'd402: toneH = `g1<<1;
		12'd403: toneH = `g1<<1;
		12'd404: toneH = `a1<<1;
		12'd405: toneH = `a1<<1;
		12'd406: toneH = `g1<<1;
		12'd407: toneH = `g1<<1;
		12'd408: toneH = `f1_u << 1;
		12'd409: toneH = `f1_u << 1;
		12'd410: toneH = `e1<<1;
		12'd411: toneH = `e1<<1;
		12'd412: toneH = `d1<<1;
		12'd413: toneH = `d1<<1;
		12'd414: toneH = `e1<<1;
		12'd415: toneH = `e1<<1;
		12'd416: toneH = `f1_u << 1;
		12'd417: toneH = `f1_u << 1;
		12'd418: toneH = `f1_u << 1;
		12'd419: toneH = `f1_u << 1;
		12'd420: toneH = `f1_u << 1;
		12'd421: toneH = `f1_u << 1;
		12'd422: toneH = `f1_u << 1;
		12'd423: toneH = `f1_u << 1;
		12'd424: toneH = `f1_u << 1;
		12'd425: toneH = `f1_u << 1;
		12'd426: toneH = `f1_u << 1;
		12'd427: toneH = `f1_u << 1;
		12'd428: toneH = `f1_u << 1;
		12'd429: toneH = `f1_u << 1;
		12'd430: toneH = `f1_u << 1;
		12'd431: toneH = `f1_u << 1;
		12'd432: toneH = `f1_u << 1;
		12'd433: toneH = `f1_u << 1;
		12'd434: toneH = `f1_u << 1;
		12'd435: toneH = `f1_u << 1;
		12'd436: toneH = `f1_u << 1;
		12'd437: toneH = `f1_u << 1;
		12'd438: toneH = `f1_u << 1;
		12'd439: toneH = `f1_u << 1;
		12'd440: toneH = `f1_u << 1;
		12'd441: toneH = `f1_u << 1;
		12'd442: toneH = `f1_u << 1;
		12'd443: toneH = `f1_u << 1;
		12'd444: toneH = `f1_u << 1;
		12'd445: toneH = `f1_u << 1;
		12'd446: toneH = `f1_u << 1;
		12'd447: toneH = `f1_u << 1;
		12'd448: toneH = `g1<<1;
		12'd449: toneH = `g1<<1;
		12'd450: toneH = `g1<<1;
		12'd451: toneH = `g1<<1;
		12'd452: toneH = `g1<<1;
		12'd453: toneH = `g1<<1;
		12'd454: toneH = `g1<<1;
		12'd455: toneH = `g1<<1;
		12'd456: toneH = `g1<<1;
		12'd457: toneH = `g1<<1;
		12'd458: toneH = `g1<<1;
		12'd459: toneH = `g1<<1;
		12'd460: toneH = `g1<<1;
		12'd461: toneH = `g1<<1;
		12'd462: toneH = `g1<<1;
		12'd463: toneH = `g1<<1;
		12'd464: toneH = `g1<<1;
		12'd465: toneH = `g1<<1;
		12'd466: toneH = `g1<<1;
		12'd467: toneH = `g1<<1;
		12'd468: toneH = `a1<<1;
		12'd469: toneH = `a1<<1;
		12'd470: toneH = `g1<<1;
		12'd471: toneH = `g1<<1;
		12'd472: toneH = `g1<<1;
		12'd473: toneH = `g1<<1;
		12'd474: toneH = `f1_u << 1;
		12'd475: toneH = `f1_u << 1;
		12'd476: toneH = `e1<<1;
		12'd477: toneH = `e1<<1;
		12'd478: toneH = `f1_u << 1;
		12'd479: toneH = `f1_u << 1;
		12'd480: toneH = `g1_u << 1;
		12'd481: toneH = `g1_u << 1;
		12'd482: toneH = `g1_u << 1;
		12'd483: toneH = `g1_u << 1;
		12'd484: toneH = `g1_u << 1;
		12'd485: toneH = `g1_u << 1;
		12'd486: toneH = `g1_u << 1;
		12'd487: toneH = `g1_u << 1;
		12'd488: toneH = `g1_u << 1;
		12'd489: toneH = `g1_u << 1;
		12'd490: toneH = `g1_u << 1;
		12'd491: toneH = `g1_u << 1;
		12'd492: toneH = `g1_u << 1;
		12'd493: toneH = `g1_u << 1;
		12'd494: toneH = `g1_u << 1;
		12'd495: toneH = `g1_u << 1;
		12'd496: toneH = `g1_u << 1;
		12'd497: toneH = `g1_u << 1;
		12'd498: toneH = `g1_u << 1;
		12'd499: toneH = `g1_u << 1;
		12'd500: toneH = `g1_u << 1;
		12'd501: toneH = `g1_u << 1;
		12'd502: toneH = `g1_u << 1;
		12'd503: toneH = `g1_u << 1;
		12'd504: toneH = `g1_u << 1;
		12'd505: toneH = `g1_u << 1;
		12'd506: toneH = `g1_u << 1;
		12'd507: toneH = `g1_u << 1;
		12'd508: toneH = `g1_u << 1;
		12'd509: toneH = `g1_u << 1;
		12'd510: toneH = `g1_u << 1;
		12'd511: toneH = `g1_u << 1;
		12'd512: toneH = `a1<<1;
		12'd513: toneH = `a1<<1;
		12'd514: toneH = `a1<<1;
		12'd515: toneH = `a1<<1;
		12'd516: toneH = `a1<<1;
		12'd517: toneH = `a1<<1;
		12'd518: toneH = `a1<<1;
		12'd519: toneH = `a1<<1;
		12'd520: toneH = `a1<<1;
		12'd521: toneH = `a1<<1;
		12'd522: toneH = `a1<<1;
		12'd523: toneH = `a1<<1;
		12'd524: toneH = `a1<<1;
		12'd525: toneH = `a1<<1;
		12'd526: toneH = `a1<<1;
		12'd527: toneH = `a1<<1;
		12'd528: toneH = `c1_u << 2;
		12'd529: toneH = `c1_u << 2;
		12'd530: toneH = `c1_u << 2;
		12'd531: toneH = `c1_u << 2;
		12'd532: toneH = `c1_u << 2;
		12'd533: toneH = `c1_u << 2;
		12'd534: toneH = `c1_u << 2;
		12'd535: toneH = `c1_u << 2;
		12'd536: toneH = `e1 << 2;
		12'd537: toneH = `e1 << 2;
		12'd538: toneH = `e1 << 2;
		12'd539: toneH = `e1 << 2;
		12'd540: toneH = `e1 << 2;
		12'd541: toneH = `e1 << 2;
		12'd542: toneH = `e1 << 2;
		12'd543: toneH = `e1 << 2;
		12'd544: toneH = `d1 << 2;
		12'd545: toneH = `d1 << 2;
		12'd546: toneH = `d1 << 2;
		12'd547: toneH = `d1 << 2;
		12'd548: toneH = `a1<<1;
		12'd549: toneH = `a1<<1;
		12'd550: toneH = `a1<<1;
		12'd551: toneH = `a1<<1;
		12'd552: toneH = `c1 << 2;
		12'd553: toneH = `c1 << 2;
		12'd554: toneH = `b1<<1;
		12'd555: toneH = `b1<<1;
		12'd556: toneH = `b1<<1;
		12'd557: toneH = `b1<<1;
		12'd558: toneH = `b1<<1;
		12'd559: toneH = `b1<<1;
		12'd560: toneH = `b1<<1;
		12'd561: toneH = `b1<<1;
		12'd562: toneH = `b1<<1;
		12'd563: toneH = `b1<<1;
		12'd564: toneH = `b1<<1;
		12'd565: toneH = `b1<<1;
		12'd566: toneH = `b1<<1;
		12'd567: toneH = `b1<<1;
		12'd568: toneH = `b1<<1;
		12'd569: toneH = `b1<<1;
		12'd570: toneH = `b1<<1;
		12'd571: toneH = `b1<<1;
		12'd572: toneH = `b1<<1;
		12'd573: toneH = `b1<<1;
		12'd574: toneH = `b1<<1;
		12'd575: toneH = `b1<<1;
		12'd576: toneH = `b1<<1;
		12'd577: toneH = `b1<<1;
		12'd578: toneH = `b1<<1;
		12'd579: toneH = `b1<<1;
		12'd580: toneH = `b1<<1;
		12'd581: toneH = `b1<<1;
		12'd582: toneH = `b1<<1;
		12'd583: toneH = `b1<<1;
		12'd584: toneH = `d1 << 2;
		12'd585: toneH = `d1 << 2;
		12'd586: toneH = `d1 << 2;
		12'd587: toneH = `d1 << 2;
		12'd588: toneH = `a1<<1;
		12'd589: toneH = `a1<<1;
		12'd590: toneH = `a1<<1;
		12'd591: toneH = `a1<<1;
		12'd592: toneH = `b1_d << 1;
		12'd593: toneH = `b1_d << 1;
		12'd594: toneH = `f1 << 2;
		12'd595: toneH = `f1 << 2;
		12'd596: toneH = `f1 << 2;
		12'd597: toneH = `f1 << 2;
		12'd598: toneH = `f1 << 2;
		12'd599: toneH = `f1 << 2;
		12'd600: toneH = `f1 << 2;
		12'd601: toneH = `f1 << 2;
		12'd602: toneH = `f1 << 2;
		12'd603: toneH = `f1 << 2;
		12'd604: toneH = `f1 << 2;
		12'd605: toneH = `f1 << 2;
		12'd606: toneH = `f1 << 2;
		12'd607: toneH = `f1 << 2;
		12'd608: toneH = `g1 << 2;
		12'd609: toneH = `g1 << 2;
		12'd610: toneH = `g1 << 2;
		12'd611: toneH = `g1 << 2;
		12'd612: toneH = `g1 << 2;
		12'd613: toneH = `g1 << 2;
		12'd614: toneH = `g1 << 2;
		12'd615: toneH = `g1 << 2;
		12'd616: toneH = `g1 << 2;
		12'd617: toneH = `g1 << 2;
		12'd618: toneH = `g1 << 2;
		12'd619: toneH = `g1 << 2;
		12'd620: toneH = `g1 << 2;
		12'd621: toneH = `g1 << 2;
		12'd622: toneH = `g1 << 2;
		12'd623: toneH = `g1 << 2;
		12'd624: toneH = `c1 << 2;
		12'd625: toneH = `c1 << 2;
		12'd626: toneH = `c1 << 2;
		12'd627: toneH = `c1 << 2;
		12'd628: toneH = `c1 << 2;
		12'd629: toneH = `c1 << 2;
		12'd630: toneH = `c1 << 2;
		12'd631: toneH = `c1 << 2;
		12'd632: toneH = `c1 << 2;
		12'd633: toneH = `c1 << 2;
		12'd634: toneH = `c1 << 2;
		12'd635: toneH = `c1 << 2;
		12'd636: toneH = `c1 << 2;
		12'd637: toneH = `c1 << 2;
		12'd638: toneH = `c1 << 2;
		12'd639: toneH = `c1 << 2;
		12'd640: toneH = `c1 << 2;
		12'd641: toneH = `c1 << 2;
		12'd642: toneH = `c1 << 2;
		12'd643: toneH = `c1 << 2;
		12'd644: toneH = `c1 << 2;
		12'd645: toneH = `c1 << 2;
		12'd646: toneH = `c1 << 2;
		12'd647: toneH = `c1 << 2;
		12'd648: toneH = `c1 << 2;
		12'd649: toneH = `c1 << 2;
		12'd650: toneH = `c1 << 2;
		12'd651: toneH = `c1 << 2;
		12'd652: toneH = `c1 << 2;
		12'd653: toneH = `c1 << 2;
		12'd654: toneH = `c1 << 2;
		12'd655: toneH = `c1 << 2;

		default : toneH = `non;
	endcase
end

always @(*) begin
	case (ibeatNum)		// 1/4 beat
		12'd0: toneM = `non;
		12'd1: toneM = `non;
		12'd2: toneM = `non;
		12'd3: toneM = `non;
		12'd4: toneM = `non;
		12'd5: toneM = `non;
		12'd6: toneM = `non;
		12'd7: toneM = `non;
		12'd8: toneM = `f1;
		12'd9: toneM = `e1;
		12'd10: toneM = `f1;
		12'd11: toneM = `e1;
		12'd12: toneM = `e1_d;
		12'd13: toneM = `e1;
		12'd14: toneM = `e1_d;
		12'd15: toneM = `d1;
		12'd16: toneM = `e1_d;
		12'd17: toneM = `d1;
		12'd18: toneM = `c1_u;
		12'd19: toneM = `d1;
		12'd20: toneM = `c1_u;
		12'd21: toneM = `c1;
		12'd22: toneM = `c1_u;
		12'd23: toneM = `c1;
		12'd24: toneM = `b1 >> 1;
		12'd25: toneM = `c1;
		12'd26: toneM = `b1 >> 1;
		12'd27: toneM = `b1_d >> 1;
		12'd28: toneM = `b1 >> 1;
		12'd29: toneM = `b1_d >> 1;
		12'd30: toneM = `a1 >> 1;
		12'd31: toneM = `b1_d >> 1;
		12'd32: toneM = `d1;
		12'd33: toneM = `d1;
		12'd34: toneM = `non;
		12'd35: toneM = `non;
		12'd36: toneM = `non;
		12'd37: toneM = `non;
		12'd38: toneM = `e1;
		12'd39: toneM = `e1;
		12'd40: toneM = `non;
		12'd41: toneM = `non;
		12'd42: toneM = `non;
		12'd43: toneM = `non;
		12'd44: toneM = `f1;
		12'd45: toneM = `f1;
		12'd46: toneM = `non;
		12'd47: toneM = `non;
		12'd48: toneM = `d1;
		12'd49: toneM = `d1;
		12'd50: toneM = `e1;
		12'd51: toneM = `e1;
		12'd52: toneM = `non;
		12'd53: toneM = `non;
		12'd54: toneM = `f1;
		12'd55: toneM = `f1;
		12'd56: toneM = `non;
		12'd57: toneM = `non;
		12'd58: toneM = `non;
		12'd59: toneM = `non;
		12'd60: toneM = `c1;
		12'd61: toneM = `c1;
		12'd62: toneM = `non;
		12'd63: toneM = `non;
		12'd64: toneM = `d1;
		12'd65: toneM = `d1;
		12'd66: toneM = `non;
		12'd67: toneM = `non;
		12'd68: toneM = `non;
		12'd69: toneM = `non;
		12'd70: toneM = `e1;
		12'd71: toneM = `e1;
		12'd72: toneM = `non;
		12'd73: toneM = `non;
		12'd74: toneM = `non;
		12'd75: toneM = `non;
		12'd76: toneM = `f1;
		12'd77: toneM = `f1;
		12'd78: toneM = `non;
		12'd79: toneM = `non;
		12'd80: toneM = `d1;
		12'd81: toneM = `d1;
		12'd82: toneM = `e1;
		12'd83: toneM = `e1;
		12'd84: toneM = `non;
		12'd85: toneM = `non;
		12'd86: toneM = `f1;
		12'd87: toneM = `f1;
		12'd88: toneM = `non;
		12'd89: toneM = `non;
		12'd90: toneM = `non;
		12'd91: toneM = `non;
		12'd92: toneM = `c1;
		12'd93: toneM = `c1;
		12'd94: toneM = `d1_d;
		12'd95: toneM = `d1_d;
		12'd96: toneM = `d1;
		12'd97: toneM = `d1;
		12'd98: toneM = `non;
		12'd99: toneM = `non;
		12'd100: toneM = `non;
		12'd101: toneM = `non;
		12'd102: toneM = `e1;
		12'd103: toneM = `e1;
		12'd104: toneM = `non;
		12'd105: toneM = `non;
		12'd106: toneM = `non;
		12'd107: toneM = `non;
		12'd108: toneM = `f1;
		12'd109: toneM = `f1;
		12'd110: toneM = `non;
		12'd111: toneM = `non;
		12'd112: toneM = `d1;
		12'd113: toneM = `d1;
		12'd114: toneM = `e1;
		12'd115: toneM = `e1;
		12'd116: toneM = `non;
		12'd117: toneM = `non;
		12'd118: toneM = `f1;
		12'd119: toneM = `f1;
		12'd120: toneM = `non;
		12'd121: toneM = `non;
		12'd122: toneM = `non;
		12'd123: toneM = `non;
		12'd124: toneM = `c1;
		12'd125: toneM = `c1;
		12'd126: toneM = `non;
		12'd127: toneM = `non;
		12'd128: toneM = `d1;
		12'd129: toneM = `d1;
		12'd130: toneM = `non;
		12'd131: toneM = `non;
		12'd132: toneM = `non;
		12'd133: toneM = `non;
		12'd134: toneM = `e1;
		12'd135: toneM = `e1;
		12'd136: toneM = `non;
		12'd137: toneM = `non;
		12'd138: toneM = `non;
		12'd139: toneM = `non;
		12'd140: toneM = `f1;
		12'd141: toneM = `f1;
		12'd142: toneM = `non;
		12'd143: toneM = `non;
		12'd144: toneM = `d1;
		12'd145: toneM = `d1;
		12'd146: toneM = `e1;
		12'd147: toneM = `e1;
		12'd148: toneM = `non;
		12'd149: toneM = `non;
		12'd150: toneM = `f1;
		12'd151: toneM = `f1;
		12'd152: toneM = `non;
		12'd153: toneM = `non;
		12'd154: toneM = `non;
		12'd155: toneM = `non;
		12'd156: toneM = `c1;
		12'd157: toneM = `c1;
		12'd158: toneM = `d1_d;
		12'd159: toneM = `d1_d;
		12'd160: toneM = `d1;
		12'd161: toneM = `d1;
		12'd162: toneM = `e1;
		12'd163: toneM = `e1;
		12'd164: toneM = `e1;
		12'd165: toneM = `e1;
		12'd166: toneM = `d1_d;
		12'd167: toneM = `d1_d;
		12'd168: toneM = `d1;
		12'd169: toneM = `d1;
		12'd170: toneM = `d1;
		12'd171: toneM = `d1;
		12'd172: toneM = `b1 >> 1;
		12'd173: toneM = `b1 >> 1;
		12'd174: toneM = `b1 >> 1;
		12'd175: toneM = `b1 >> 1;
		12'd176: toneM = `g1_d >> 1;
		12'd177: toneM = `g1_d >> 1;
		12'd178: toneM = `g1_d >> 1;
		12'd179: toneM = `g1_d >> 1;
		12'd180: toneM = `e1;
		12'd181: toneM = `e1;
		12'd182: toneM = `d1;
		12'd183: toneM = `d1;
		12'd184: toneM = `d1;
		12'd185: toneM = `d1;
		12'd186: toneM = `d1_d;
		12'd187: toneM = `d1_d;
		12'd188: toneM = `d1;
		12'd189: toneM = `d1;
		12'd190: toneM = `e1;
		12'd191: toneM = `e1;
		12'd192: toneM = `f1;
		12'd193: toneM = `f1;
		12'd194: toneM = `f1;
		12'd195: toneM = `f1;
		12'd196: toneM = `f1;
		12'd197: toneM = `f1;
		12'd198: toneM = `f1;
		12'd199: toneM = `f1;
		12'd200: toneM = `c1;
		12'd201: toneM = `d1_d;
		12'd202: toneM = `d1;
		12'd203: toneM = `e1_d;
		12'd204: toneM = `e1;
		12'd205: toneM = `e1_d;
		12'd206: toneM = `d1;
		12'd207: toneM = `c1;
		12'd208: toneM = `c1;
		12'd209: toneM = `d1_d;
		12'd210: toneM = `d1;
		12'd211: toneM = `e1_d;
		12'd212: toneM = `e1;
		12'd213: toneM = `f1;
		12'd214: toneM = `f1_u;
		12'd215: toneM = `g1;
		12'd216: toneM = `g1_u;
		12'd217: toneM = `g1;
		12'd218: toneM = `f1_u;
		12'd219: toneM = `f1;
		12'd220: toneM = `e1;
		12'd221: toneM = `d1_u;
		12'd222: toneM = `d1;
		12'd223: toneM = `c1;
		12'd224: toneM = `d1;
		12'd225: toneM = `d1;
		12'd226: toneM = `e1;
		12'd227: toneM = `e1;
		12'd228: toneM = `e1;
		12'd229: toneM = `e1;
		12'd230: toneM = `d1_d;
		12'd231: toneM = `d1_d;
		12'd232: toneM = `d1;
		12'd233: toneM = `d1;
		12'd234: toneM = `d1;
		12'd235: toneM = `d1;
		12'd236: toneM = `b1 >> 1;
		12'd237: toneM = `b1 >> 1;
		12'd238: toneM = `b1 >> 1;
		12'd239: toneM = `b1 >> 1;
		12'd240: toneM = `g1_d >> 1;
		12'd241: toneM = `g1_d >> 1;
		12'd242: toneM = `g1_d >> 1;
		12'd243: toneM = `g1_d >> 1;
		12'd244: toneM = `e1;
		12'd245: toneM = `e1;
		12'd246: toneM = `d1;
		12'd247: toneM = `d1;
		12'd248: toneM = `d1;
		12'd249: toneM = `d1;
		12'd250: toneM = `c1_u;
		12'd251: toneM = `c1_u;
		12'd252: toneM = `b1 >> 1;
		12'd253: toneM = `b1 >> 1;
		12'd254: toneM = `d1_d;
		12'd255: toneM = `d1_d;
		12'd256: toneM = `d1;
		12'd257: toneM = `d1;
		12'd258: toneM = `d1;
		12'd259: toneM = `d1;
		12'd260: toneM = `d1;
		12'd261: toneM = `d1;
		12'd262: toneM = `d1;
		12'd263: toneM = `d1;
		12'd264: toneM = `c1_u;
		12'd265: toneM = `c1_u;
		12'd266: toneM = `c1_u;
		12'd267: toneM = `c1_u;
		12'd268: toneM = `c1_u;
		12'd269: toneM = `c1_u;
		12'd270: toneM = `c1_u;
		12'd271: toneM = `c1_u;
		12'd272: toneM = `b1 >> 1;
		12'd273: toneM = `b1 >> 1;
		12'd274: toneM = `b1 >> 1;
		12'd275: toneM = `b1 >> 1;
		12'd276: toneM = `b1 >> 1;
		12'd277: toneM = `b1 >> 1;
		12'd278: toneM = `b1 >> 1;
		12'd279: toneM = `b1 >> 1;
		12'd280: toneM = `c1_u;
		12'd281: toneM = `c1_u;
		12'd282: toneM = `c1_u;
		12'd283: toneM = `c1_u;
		12'd284: toneM = `c1_u;
		12'd285: toneM = `c1_u;
		12'd286: toneM = `c1_u;
		12'd287: toneM = `c1_u;
		12'd288: toneM = `d1;
		12'd289: toneM = `d1;
		12'd290: toneM = `c1_u;
		12'd291: toneM = `c1_u;
		12'd292: toneM = `b1 >> 1;
		12'd293: toneM = `b1 >> 1;
		12'd294: toneM = `a1 >> 1;
		12'd295: toneM = `a1 >> 1;
		12'd296: toneM = `g1 >> 1;
		12'd297: toneM = `g1 >> 1;
		12'd298: toneM = `g1 >> 1;
		12'd299: toneM = `g1 >> 1;
		12'd300: toneM = `d1;
		12'd301: toneM = `d1;
		12'd302: toneM = `c1;
		12'd303: toneM = `c1;
		12'd304: toneM = `b1 >> 1;
		12'd305: toneM = `b1 >> 1;
		12'd306: toneM = `a1 >> 1;
		12'd307: toneM = `a1 >> 1;
		12'd308: toneM = `g1 >> 1;
		12'd309: toneM = `g1 >> 1;
		12'd310: toneM = `g1 >> 1;
		12'd311: toneM = `g1 >> 1;
		12'd312: toneM = `d1;
		12'd313: toneM = `d1;
		12'd314: toneM = `c1_u;
		12'd315: toneM = `c1_u;
		12'd316: toneM = `b1 >> 1;
		12'd317: toneM = `b1 >> 1;
		12'd318: toneM = `c1_u;
		12'd319: toneM = `c1_u;
		12'd320: toneM = `e1;
		12'd321: toneM = `e1;
		12'd322: toneM = `e1;
		12'd323: toneM = `e1;
		12'd324: toneM = `g1 >> 1;
		12'd325: toneM = `a1 >> 1;
		12'd326: toneM = `b1 >> 1;
		12'd327: toneM = `c1_u;
		12'd328: toneM = `d1;
		12'd329: toneM = `d1;
		12'd330: toneM = `d1;
		12'd331: toneM = `d1;
		12'd332: toneM = `f1_u >> 1;
		12'd333: toneM = `g1 >> 1;
		12'd334: toneM = `a1 >> 1;
		12'd335: toneM = `b1 >> 1;
		12'd336: toneM = `c1_u;
		12'd337: toneM = `c1_u;
		12'd338: toneM = `c1_u;
		12'd339: toneM = `c1_u;
		12'd340: toneM = `g1 >> 1;
		12'd341: toneM = `a1 >> 1;
		12'd342: toneM = `b1 >> 1;
		12'd343: toneM = `c1;
		12'd344: toneM = `d1;
		12'd345: toneM = `d1;
		12'd346: toneM = `d1;
		12'd347: toneM = `d1;
		12'd348: toneM = `f1_u >> 1;
		12'd349: toneM = `g1 >> 1;
		12'd350: toneM = `a1 >> 1;
		12'd351: toneM = `b1 >> 1;
		12'd352: toneM = `d1;
		12'd353: toneM = `d1;
		12'd354: toneM = `c1_u;
		12'd355: toneM = `c1_u;
		12'd356: toneM = `b1 >> 1;
		12'd357: toneM = `b1 >> 1;
		12'd358: toneM = `a1 >> 1;
		12'd359: toneM = `a1 >> 1;
		12'd360: toneM = `g1 >> 1;
		12'd361: toneM = `g1 >> 1;
		12'd362: toneM = `g1 >> 1;
		12'd363: toneM = `g1 >> 1;
		12'd364: toneM = `d1;
		12'd365: toneM = `d1;
		12'd366: toneM = `c1_u;
		12'd367: toneM = `c1_u;
		12'd368: toneM = `b1 >> 1;
		12'd369: toneM = `b1 >> 1;
		12'd370: toneM = `a1 >> 1;
		12'd371: toneM = `a1 >> 1;
		12'd372: toneM = `b1 >> 1;
		12'd373: toneM = `b1 >> 1;
		12'd374: toneM = `g1 >> 1;
		12'd375: toneM = `g1 >> 1;
		12'd376: toneM = `d1;
		12'd377: toneM = `d1;
		12'd378: toneM = `e1;
		12'd379: toneM = `e1;
		12'd380: toneM = `f1_u;
		12'd381: toneM = `f1_u;
		12'd382: toneM = `g1;
		12'd383: toneM = `g1;
		12'd384: toneM = `a1;
		12'd385: toneM = `a1;
		12'd386: toneM = `b1;
		12'd387: toneM = `b1;
		12'd388: toneM = `a1;
		12'd389: toneM = `a1;
		12'd390: toneM = `g1;
		12'd391: toneM = `g1;
		12'd392: toneM = `a1;
		12'd393: toneM = `a1;
		12'd394: toneM = `non;
		12'd395: toneM = `non;
		12'd396: toneM = `a1;
		12'd397: toneM = `a1;
		12'd398: toneM = `b1;
		12'd399: toneM = `b1;
		12'd400: toneM = `a1;
		12'd401: toneM = `a1;
		12'd402: toneM = `g1;
		12'd403: toneM = `g1;
		12'd404: toneM = `f1_u;
		12'd405: toneM = `f1_u;
		12'd406: toneM = `g1;
		12'd407: toneM = `g1;
		12'd408: toneM = `a1;
		12'd409: toneM = `a1;
		12'd410: toneM = `e1;
		12'd411: toneM = `e1;
		12'd412: toneM = `g1;
		12'd413: toneM = `g1;
		12'd414: toneM = `f1_u;
		12'd415: toneM = `f1_u;
		12'd416: toneM = `b1 >> 1;
		12'd417: toneM = `c1;
		12'd418: toneM = `d1_d;
		12'd419: toneM = `d1;
		12'd420: toneM = `d1_u;
		12'd421: toneM = `e1;
		12'd422: toneM = `f1;
		12'd423: toneM = `g1_d;
		12'd424: toneM = `g1;
		12'd425: toneM = `g1_u;
		12'd426: toneM = `a1;
		12'd427: toneM = `a1_u;
		12'd428: toneM = `b1;
		12'd429: toneM = `c1 << 1;
		12'd430: toneM = `c1_u << 1;
		12'd431: toneM = `d1 << 1;
		12'd432: toneM = `d1_u << 1;
		12'd433: toneM = `d1 << 1;
		12'd434: toneM = `d1_d << 1;
		12'd435: toneM = `c1 << 1;
		12'd436: toneM = `b1;
		12'd437: toneM = `b1_d;
		12'd438: toneM = `a1;
		12'd439: toneM = `a1_d;
		12'd440: toneM = `g1;
		12'd441: toneM = `g1_d;
		12'd442: toneM = `f1;
		12'd443: toneM = `e1;
		12'd444: toneM = `e1_d;
		12'd445: toneM = `d1;
		12'd446: toneM = `d1_d;
		12'd447: toneM = `c1;
		12'd448: toneM = `c1;
		12'd449: toneM = `c1_u;
		12'd450: toneM = `d1;
		12'd451: toneM = `d1_u;
		12'd452: toneM = `e1;
		12'd453: toneM = `f1;
		12'd454: toneM = `f1_u;
		12'd455: toneM = `g1;
		12'd456: toneM = `g1_u;
		12'd457: toneM = `a1;
		12'd458: toneM = `b1_d;
		12'd459: toneM = `b1;
		12'd460: toneM = `c1 << 1;
		12'd461: toneM = `c1_u << 1;
		12'd462: toneM = `d1 << 1;
		12'd463: toneM = `d1_u << 1;
		12'd464: toneM = `e1 << 1;
		12'd465: toneM = `e1_d << 1;
		12'd466: toneM = `d1 << 1;
		12'd467: toneM = `d1_d << 1;
		12'd468: toneM = `c1_u << 1;
		12'd469: toneM = `b1;
		12'd470: toneM = `b1_d;
		12'd471: toneM = `a1;
		12'd472: toneM = `a1_d;
		12'd473: toneM = `g1;
		12'd474: toneM = `g1_d;
		12'd475: toneM = `f1;
		12'd476: toneM = `e1;
		12'd477: toneM = `e1_d;
		12'd478: toneM = `d1;
		12'd479: toneM = `d1_d;
		12'd480: toneM = `d1_d;
		12'd481: toneM = `d1;
		12'd482: toneM = `d1_u;
		12'd483: toneM = `e1;
		12'd484: toneM = `f1;
		12'd485: toneM = `f1_u;
		12'd486: toneM = `g1;
		12'd487: toneM = `g1_u;
		12'd488: toneM = `a1;
		12'd489: toneM = `a1_u;
		12'd490: toneM = `b1;
		12'd491: toneM = `c1 << 1;
		12'd492: toneM = `c1_u << 1;
		12'd493: toneM = `d1 << 1;
		12'd494: toneM = `d1_u << 1;
		12'd495: toneM = `e1 << 1;
		12'd496: toneM = `f1 << 1;
		12'd497: toneM = `e1 << 1;
		12'd498: toneM = `e1_d << 1;
		12'd499: toneM = `d1 << 1;
		12'd500: toneM = `d1_d << 1;
		12'd501: toneM = `c1 << 1;
		12'd502: toneM = `b1;
		12'd503: toneM = `b1_d;
		12'd504: toneM = `a1;
		12'd505: toneM = `a1_d;
		12'd506: toneM = `g1;
		12'd507: toneM = `g1_d;
		12'd508: toneM = `f1;
		12'd509: toneM = `e1;
		12'd510: toneM = `e1_d;
		12'd511: toneM = `d1;
		12'd512: toneM = `d1;
		12'd513: toneM = `d1_u;
		12'd514: toneM = `e1;
		12'd515: toneM = `f1;
		12'd516: toneM = `f1_u;
		12'd517: toneM = `g1;
		12'd518: toneM = `g1_u;
		12'd519: toneM = `a1;
		12'd520: toneM = `a1_u;
		12'd521: toneM = `b1;
		12'd522: toneM = `c1 << 1;
		12'd523: toneM = `c1_u << 1;
		12'd524: toneM = `d1 << 1;
		12'd525: toneM = `d1_u << 1;
		12'd526: toneM = `e1 << 1;
		12'd527: toneM = `f1 << 1;
		12'd528: toneM = `f1_u << 1;
		12'd529: toneM = `f1 << 1;
		12'd530: toneM = `e1 << 1;
		12'd531: toneM = `e1_d << 1;
		12'd532: toneM = `d1 << 1;
		12'd533: toneM = `c1_u << 1;
		12'd534: toneM = `c1 << 1;
		12'd535: toneM = `b1;
		12'd536: toneM = `b1_d;
		12'd537: toneM = `a1;
		12'd538: toneM = `a1_d;
		12'd539: toneM = `g1;
		12'd540: toneM = `g1_d;
		12'd541: toneM = `f1;
		12'd542: toneM = `e1;
		12'd543: toneM = `e1_d;
		12'd544: toneM = `a1;
		12'd545: toneM = `a1;
		12'd546: toneM = `a1;
		12'd547: toneM = `a1;
		12'd548: toneM = `d1 << 1;
		12'd549: toneM = `d1 << 1;
		12'd550: toneM = `d1 << 1;
		12'd551: toneM = `d1 << 1;
		12'd552: toneM = `a1;
		12'd553: toneM = `a1;
		12'd554: toneM = `d1;
		12'd555: toneM = `e1;
		12'd556: toneM = `f1_u;
		12'd557: toneM = `g1;
		12'd558: toneM = `g1_u;
		12'd559: toneM = `a1_u;
		12'd560: toneM = `b1;
		12'd561: toneM = `b1;
		12'd562: toneM = `c1 << 1;
		12'd563: toneM = `c1 << 1;
		12'd564: toneM = `a1;
		12'd565: toneM = `a1;
		12'd566: toneM = `c1 << 1;
		12'd567: toneM = `c1 << 1;
		12'd568: toneM = `g1;
		12'd569: toneM = `g1;
		12'd570: toneM = `b1;
		12'd571: toneM = `b1;
		12'd572: toneM = `f1;
		12'd573: toneM = `f1;
		12'd574: toneM = `g1;
		12'd575: toneM = `g1;
		12'd576: toneM = `a1;
		12'd577: toneM = `a1;
		12'd578: toneM = `c1 << 1;
		12'd579: toneM = `c1 << 1;
		12'd580: toneM = `d1 << 1;
		12'd581: toneM = `d1 << 1;
		12'd582: toneM = `non;
		12'd583: toneM = `non;
		12'd584: toneM = `a1;
		12'd585: toneM = `a1;
		12'd586: toneM = `a1;
		12'd587: toneM = `a1;
		12'd588: toneM = `c1 << 1;
		12'd589: toneM = `c1 << 1;
		12'd590: toneM = `c1 << 1;
		12'd591: toneM = `c1 << 1;
		12'd592: toneM = `d1 << 1;
		12'd593: toneM = `d1 << 1;
		12'd594: toneM = `f1;
		12'd595: toneM = `g1;
		12'd596: toneM = `a1;
		12'd597: toneM = `b1;
		12'd598: toneM = `c1 << 1;
		12'd599: toneM = `d1 << 1;
		12'd600: toneM = `e1 << 1;
		12'd601: toneM = `e1 << 1;
		12'd602: toneM = `f1 << 1;
		12'd603: toneM = `f1 << 1;
		12'd604: toneM = `d1 << 1;
		12'd605: toneM = `d1 << 1;
		12'd606: toneM = `f1 << 1;
		12'd607: toneM = `f1 << 1;
		12'd608: toneM = `d1 << 1;
		12'd609: toneM = `d1 << 1;
		12'd610: toneM = `f1 << 1;
		12'd611: toneM = `f1 << 1;
		12'd612: toneM = `d1 << 1;
		12'd613: toneM = `d1 << 1;
		12'd614: toneM = `f1 << 1;
		12'd615: toneM = `f1 << 1;
		12'd616: toneM = `d1 << 1;
		12'd617: toneM = `d1 << 1;
		12'd618: toneM = `f1 << 1;
		12'd619: toneM = `f1 << 1;
		12'd620: toneM = `d1 << 1;
		12'd621: toneM = `d1 << 1;
		12'd622: toneM = `f1 << 1;
		12'd623: toneM = `f1 << 1;
		12'd624: toneM = `e1 << 1;
		12'd625: toneM = `e1 << 1;
		12'd626: toneM = `f1 << 1;
		12'd627: toneM = `f1 << 1;
		12'd628: toneM = `e1 << 1;
		12'd629: toneM = `e1 << 1;
		12'd630: toneM = `f1 << 1;
		12'd631: toneM = `f1 << 1;
		12'd632: toneM = `e1 << 1;
		12'd633: toneM = `e1 << 1;
		12'd634: toneM = `f1 << 1;
		12'd635: toneM = `f1 << 1;
		12'd636: toneM = `e1 << 1;
		12'd637: toneM = `e1 << 1;
		12'd638: toneM = `f1 << 1;
		12'd639: toneM = `f1 << 1;
		12'd640: toneM = `e1 << 1;
		12'd641: toneM = `e1 << 1;
		12'd642: toneM = `f1 << 1;
		12'd643: toneM = `f1 << 1;
		12'd644: toneM = `e1 << 1;
		12'd645: toneM = `e1 << 1;
		12'd646: toneM = `f1 << 1;
		12'd647: toneM = `f1 << 1;
		12'd648: toneM = `e1 << 1;
		12'd649: toneM = `e1 << 1;
		12'd650: toneM = `f1 << 1;
		12'd651: toneM = `f1 << 1;
		12'd652: toneM = `e1 << 1;
		12'd653: toneM = `e1 << 1;
		12'd654: toneM = `b1;
		12'd655: toneM = `b1;


		default : toneM = `non;
	endcase
end

always @(*) begin
	case (ibeatNum)		// 1/4 beat
		12'd0: toneL = `b1 >> 1;
		12'd1: toneL = `b1_d >> 1;
		12'd2: toneL = `a1 >> 1;
		12'd3: toneL = `a1_d >> 1;
		12'd4: toneL = `a1 >> 1;
		12'd5: toneL = `g1_u >> 1;
		12'd6: toneL = `g1 >> 1;
		12'd7: toneL = `f1_u >> 1;
		12'd8: toneL = `g1 >> 1;
		12'd9: toneL = `g1_d >> 1;
		12'd10: toneL = `f1 >> 1;
		12'd11: toneL = `e1 >> 1;
		12'd12: toneL = `f1 >> 1;
		12'd13: toneL = `e1 >> 1;
		12'd14: toneL = `d1_u >> 1;
		12'd15: toneL = `d1 >> 1;
		12'd16: toneL = `e1_d >> 1;
		12'd17: toneL = `d1 >> 1;
		12'd18: toneL = `c1_u >> 1;
		12'd19: toneL = `c1_u >> 1;
		12'd20: toneL = `d1_d >> 1;
		12'd21: toneL = `c1_u >> 1;
		12'd22: toneL = `b1 >> 2;
		12'd23: toneL = `a1_u >> 2;
		12'd24: toneL = `b1 >> 2;
		12'd25: toneL = `a1_u >> 2;
		12'd26: toneL = `a1 >> 2;
		12'd27: toneL = `g1_u >> 2;
		12'd28: toneL = `a1 >> 2;
		12'd29: toneL = `g1_u >> 2;
		12'd30: toneL = `g1 >> 2;
		12'd31: toneL = `g1_d >> 2;
		12'd32: toneL = `b1 >> 2;
		12'd33: toneL = `b1 >> 2;
		12'd34: toneL = `b1 >> 2;
		12'd35: toneL = `b1 >> 2;
		12'd36: toneL = `d1 >> 1;
		12'd37: toneL = `d1 >> 1;
		12'd38: toneL = `e1 >> 1;
		12'd39: toneL = `e1 >> 1;
		12'd40: toneL = `b1 >> 2;
		12'd41: toneL = `b1 >> 2;
		12'd42: toneL = `f1 >> 1;
		12'd43: toneL = `f1 >> 1;
		12'd44: toneL = `e1 >> 1;
		12'd45: toneL = `e1 >> 1;
		12'd46: toneL = `d1 >> 1;
		12'd47: toneL = `d1 >> 1;
		12'd48: toneL = `b1 >> 2;
		12'd49: toneL = `b1 >> 2;
		12'd50: toneL = `b1 >> 2;
		12'd51: toneL = `b1 >> 2;
		12'd52: toneL = `d1 >> 1;
		12'd53: toneL = `d1 >> 1;
		12'd54: toneL = `e1 >> 1;
		12'd55: toneL = `e1 >> 1;
		12'd56: toneL = `b1 >> 2;
		12'd57: toneL = `b1 >> 2;
		12'd58: toneL = `d1 >> 1;
		12'd59: toneL = `d1 >> 1;
		12'd60: toneL = `a1_u >> 2;
		12'd61: toneL = `a1_u >> 2;
		12'd62: toneL = `c1 >> 1;
		12'd63: toneL = `c1 >> 1;
		12'd64: toneL = `b1 >> 2;
		12'd65: toneL = `b1 >> 2;
		12'd66: toneL = `b1 >> 2;
		12'd67: toneL = `b1 >> 2;
		12'd68: toneL = `d1 >> 1;
		12'd69: toneL = `d1 >> 1;
		12'd70: toneL = `e1 >> 1;
		12'd71: toneL = `e1 >> 1;
		12'd72: toneL = `b1 >> 2;
		12'd73: toneL = `b1 >> 2;
		12'd74: toneL = `f1 >> 1;
		12'd75: toneL = `f1 >> 1;
		12'd76: toneL = `e1 >> 1;
		12'd77: toneL = `e1 >> 1;
		12'd78: toneL = `d1 >> 1;
		12'd79: toneL = `d1 >> 1;
		12'd80: toneL = `b1 >> 2;
		12'd81: toneL = `b1 >> 2;
		12'd82: toneL = `b1 >> 2;
		12'd83: toneL = `b1 >> 2;
		12'd84: toneL = `d1 >> 1;
		12'd85: toneL = `d1 >> 1;
		12'd86: toneL = `e1 >> 1;
		12'd87: toneL = `e1 >> 1;
		12'd88: toneL = `b1 >> 2;
		12'd89: toneL = `b1 >> 2;
		12'd90: toneL = `d1 >> 1;
		12'd91: toneL = `d1 >> 1;
		12'd92: toneL = `a1_u >> 2;
		12'd93: toneL = `a1_u >> 2;
		12'd94: toneL = `c1 >> 1;
		12'd95: toneL = `c1 >> 1;
		12'd96: toneL = `b1 >> 2;
		12'd97: toneL = `b1 >> 2;
		12'd98: toneL = `b1 >> 2;
		12'd99: toneL = `b1 >> 2;
		12'd100: toneL = `d1 >> 1;
		12'd101: toneL = `d1 >> 1;
		12'd102: toneL = `e1 >> 1;
		12'd103: toneL = `e1 >> 1;
		12'd104: toneL = `b1 >> 2;
		12'd105: toneL = `b1 >> 2;
		12'd106: toneL = `f1 >> 1;
		12'd107: toneL = `f1 >> 1;
		12'd108: toneL = `e1 >> 1;
		12'd109: toneL = `e1 >> 1;
		12'd110: toneL = `d1 >> 1;
		12'd111: toneL = `d1 >> 1;
		12'd112: toneL = `b1 >> 2;
		12'd113: toneL = `b1 >> 2;
		12'd114: toneL = `b1 >> 2;
		12'd115: toneL = `b1 >> 2;
		12'd116: toneL = `d1 >> 1;
		12'd117: toneL = `d1 >> 1;
		12'd118: toneL = `e1 >> 1;
		12'd119: toneL = `e1 >> 1;
		12'd120: toneL = `b1 >> 2;
		12'd121: toneL = `b1 >> 2;
		12'd122: toneL = `d1 >> 1;
		12'd123: toneL = `d1 >> 1;
		12'd124: toneL = `a1_u >> 2;
		12'd125: toneL = `a1_u >> 2;
		12'd126: toneL = `c1 >> 1;
		12'd127: toneL = `c1 >> 1;
		12'd128: toneL = `b1 >> 2;
		12'd129: toneL = `b1 >> 2;
		12'd130: toneL = `b1 >> 2;
		12'd131: toneL = `b1 >> 2;
		12'd132: toneL = `d1 >> 1;
		12'd133: toneL = `d1 >> 1;
		12'd134: toneL = `e1 >> 1;
		12'd135: toneL = `e1 >> 1;
		12'd136: toneL = `b1 >> 2;
		12'd137: toneL = `b1 >> 2;
		12'd138: toneL = `f1 >> 1;
		12'd139: toneL = `f1 >> 1;
		12'd140: toneL = `e1 >> 1;
		12'd141: toneL = `e1 >> 1;
		12'd142: toneL = `d1 >> 1;
		12'd143: toneL = `d1 >> 1;
		12'd144: toneL = `b1 >> 2;
		12'd145: toneL = `b1 >> 2;
		12'd146: toneL = `b1 >> 2;
		12'd147: toneL = `b1 >> 2;
		12'd148: toneL = `d1 >> 1;
		12'd149: toneL = `d1 >> 1;
		12'd150: toneL = `e1 >> 1;
		12'd151: toneL = `e1 >> 1;
		12'd152: toneL = `b1 >> 2;
		12'd153: toneL = `b1 >> 2;
		12'd154: toneL = `d1 >> 1;
		12'd155: toneL = `d1 >> 1;
		12'd156: toneL = `a1_u >> 2;
		12'd157: toneL = `a1_u >> 2;
		12'd158: toneL = `c1 >> 1;
		12'd159: toneL = `c1 >> 1;
		12'd160: toneL = `b1 >> 2;
		12'd161: toneL = `b1 >> 2;
		12'd162: toneL = `f1_u >> 1;
		12'd163: toneL = `f1_u >> 1;
		12'd164: toneL = `b1 >> 2;
		12'd165: toneL = `b1 >> 2;
		12'd166: toneL = `f1_u >> 1;
		12'd167: toneL = `f1_u >> 1;
		12'd168: toneL = `b1 >> 2;
		12'd169: toneL = `b1 >> 2;
		12'd170: toneL = `f1_u >> 1;
		12'd171: toneL = `f1_u >> 1;
		12'd172: toneL = `b1 >> 2;
		12'd173: toneL = `b1 >> 2;
		12'd174: toneL = `f1_u >> 1;
		12'd175: toneL = `f1_u >> 1;
		12'd176: toneL = `b1 >> 2;
		12'd177: toneL = `b1 >> 2;
		12'd178: toneL = `f1_u >> 1;
		12'd179: toneL = `f1_u >> 1;
		12'd180: toneL = `b1 >> 2;
		12'd181: toneL = `b1 >> 2;
		12'd182: toneL = `f1_u >> 1;
		12'd183: toneL = `f1_u >> 1;
		12'd184: toneL = `b1 >> 2;
		12'd185: toneL = `b1 >> 2;
		12'd186: toneL = `f1_u >> 1;
		12'd187: toneL = `f1_u >> 1;
		12'd188: toneL = `b1 >> 2;
		12'd189: toneL = `b1 >> 2;
		12'd190: toneL = `f1 >> 1;
		12'd191: toneL = `f1 >> 1;
		12'd192: toneL = `b1 >> 2;
		12'd193: toneL = `b1 >> 2;
		12'd194: toneL = `g1 >> 1;
		12'd195: toneL = `g1 >> 1;
		12'd196: toneL = `c1 >> 1;
		12'd197: toneL = `c1 >> 1;
		12'd198: toneL = `g1 >> 1;
		12'd199: toneL = `g1 >> 1;
		12'd200: toneL = `c1 >> 1;
		12'd201: toneL = `c1 >> 1;
		12'd202: toneL = `g1 >> 1;
		12'd203: toneL = `g1 >> 1;
		12'd204: toneL = `c1 >> 1;
		12'd205: toneL = `c1 >> 1;
		12'd206: toneL = `g1 >> 1;
		12'd207: toneL = `g1 >> 1;
		12'd208: toneL = `c1 >> 1;
		12'd209: toneL = `c1 >> 1;
		12'd210: toneL = `g1 >> 1;
		12'd211: toneL = `g1 >> 1;
		12'd212: toneL = `a1 >> 1;
		12'd213: toneL = `a1 >> 1;
		12'd214: toneL = `g1 >> 1;
		12'd215: toneL = `g1 >> 1;
		12'd216: toneL = `f1_u >> 1;
		12'd217: toneL = `f1_u >> 1;
		12'd218: toneL = `e1 >> 1;
		12'd219: toneL = `e1 >> 1;
		12'd220: toneL = `d1 >> 1;
		12'd221: toneL = `d1 >> 1;
		12'd222: toneL = `c1 >> 1;
		12'd223: toneL = `c1 >> 1;
		12'd224: toneL = `b1 >> 2;
		12'd225: toneL = `b1 >> 2;
		12'd226: toneL = `f1 >> 1;
		12'd227: toneL = `f1 >> 1;
		12'd228: toneL = `b1 >> 2;
		12'd229: toneL = `b1 >> 2;
		12'd230: toneL = `f1_u >> 1;
		12'd231: toneL = `f1_u >> 1;
		12'd232: toneL = `b1 >> 2;
		12'd233: toneL = `b1 >> 2;
		12'd234: toneL = `f1_u >> 1;
		12'd235: toneL = `f1_u >> 1;
		12'd236: toneL = `b1 >> 2;
		12'd237: toneL = `b1 >> 2;
		12'd238: toneL = `f1_u >> 1;
		12'd239: toneL = `f1_u >> 1;
		12'd240: toneL = `b1 >> 2;
		12'd241: toneL = `b1 >> 2;
		12'd242: toneL = `f1_u >> 1;
		12'd243: toneL = `f1_u >> 1;
		12'd244: toneL = `b1 >> 2;
		12'd245: toneL = `b1 >> 2;
		12'd246: toneL = `f1_u >> 1;
		12'd247: toneL = `f1_u >> 1;
		12'd248: toneL = `b1 >> 2;
		12'd249: toneL = `b1 >> 2;
		12'd250: toneL = `f1_u >> 1;
		12'd251: toneL = `f1_u >> 1;
		12'd252: toneL = `b1 >> 2;
		12'd253: toneL = `b1 >> 2;
		12'd254: toneL = `f1 >> 1;
		12'd255: toneL = `f1 >> 1;
		12'd256: toneL = `a1 >> 2;
		12'd257: toneL = `a1 >> 2;
		12'd258: toneL = `e1_d >> 1;
		12'd259: toneL = `e1_d >> 1;
		12'd260: toneL = `a1 >> 2;
		12'd261: toneL = `a1 >> 2;
		12'd262: toneL = `e1 >> 1;
		12'd263: toneL = `e1 >> 1;
		12'd264: toneL = `a1 >> 2;
		12'd265: toneL = `a1 >> 2;
		12'd266: toneL = `e1 >> 1;
		12'd267: toneL = `e1 >> 1;
		12'd268: toneL = `a1 >> 2;
		12'd269: toneL = `a1 >> 2;
		12'd270: toneL = `e1 >> 1;
		12'd271: toneL = `e1 >> 1;
		12'd272: toneL = `a1 >> 2;
		12'd273: toneL = `a1 >> 2;
		12'd274: toneL = `e1 >> 1;
		12'd275: toneL = `e1 >> 1;
		12'd276: toneL = `d1 >> 1;
		12'd277: toneL = `d1 >> 1;
		12'd278: toneL = `c1_u >> 1;
		12'd279: toneL = `c1_u >> 1;
		12'd280: toneL = `d1 >> 1;
		12'd281: toneL = `d1 >> 1;
		12'd282: toneL = `c1_u >> 1;
		12'd283: toneL = `c1_u >> 1;
		12'd284: toneL = `a1 >> 2;
		12'd285: toneL = `a1 >> 2;
		12'd286: toneL = `g1_u >> 2;
		12'd287: toneL = `g1_u >> 2;
		12'd288: toneL = `g1 >> 2;
		12'd289: toneL = `g1 >> 2;
		12'd290: toneL = `c1_u >> 1;
		12'd291: toneL = `c1_u >> 1;
		12'd292: toneL = `g1 >> 2;
		12'd293: toneL = `g1 >> 2;
		12'd294: toneL = `d1 >> 1;
		12'd295: toneL = `d1 >> 1;
		12'd296: toneL = `g1 >> 2;
		12'd297: toneL = `g1 >> 2;
		12'd298: toneL = `d1 >> 1;
		12'd299: toneL = `d1 >> 1;
		12'd300: toneL = `g1 >> 2;
		12'd301: toneL = `g1 >> 2;
		12'd302: toneL = `d1 >> 1;
		12'd303: toneL = `d1 >> 1;
		12'd304: toneL = `g1 >> 2;
		12'd305: toneL = `g1 >> 2;
		12'd306: toneL = `d1 >> 1;
		12'd307: toneL = `d1 >> 1;
		12'd308: toneL = `g1 >> 2;
		12'd309: toneL = `g1 >> 2;
		12'd310: toneL = `d1 >> 1;
		12'd311: toneL = `d1 >> 1;
		12'd312: toneL = `g1 >> 2;
		12'd313: toneL = `g1 >> 2;
		12'd314: toneL = `d1 >> 1;
		12'd315: toneL = `d1 >> 1;
		12'd316: toneL = `g1 >> 2;
		12'd317: toneL = `g1 >> 2;
		12'd318: toneL = `a1_d >> 2;
		12'd319: toneL = `a1_d >> 2;
		12'd320: toneL = `a1 >> 2;
		12'd321: toneL = `a1 >> 2;
		12'd322: toneL = `e1 >> 1;
		12'd323: toneL = `e1 >> 1;
		12'd324: toneL = `a1 >> 2;
		12'd325: toneL = `a1 >> 2;
		12'd326: toneL = `e1 >> 1;
		12'd327: toneL = `e1 >> 1;
		12'd328: toneL = `a1 >> 2;
		12'd329: toneL = `a1 >> 2;
		12'd330: toneL = `e1 >> 1;
		12'd331: toneL = `e1 >> 1;
		12'd332: toneL = `a1 >> 2;
		12'd333: toneL = `a1 >> 2;
		12'd334: toneL = `e1 >> 1;
		12'd335: toneL = `e1 >> 1;
		12'd336: toneL = `a1 >> 2;
		12'd337: toneL = `a1 >> 2;
		12'd338: toneL = `e1 >> 1;
		12'd339: toneL = `e1 >> 1;
		12'd340: toneL = `a1 >> 2;
		12'd341: toneL = `a1 >> 2;
		12'd342: toneL = `e1 >> 1;
		12'd343: toneL = `e1 >> 1;
		12'd344: toneL = `a1 >> 2;
		12'd345: toneL = `a1 >> 2;
		12'd346: toneL = `e1 >> 1;
		12'd347: toneL = `e1 >> 1;
		12'd348: toneL = `a1 >> 2;
		12'd349: toneL = `a1 >> 2;
		12'd350: toneL = `e1 >> 1;
		12'd351: toneL = `e1 >> 1;
		12'd352: toneL = `g1 >> 2;
		12'd353: toneL = `g1 >> 2;
		12'd354: toneL = `d1 >> 1;
		12'd355: toneL = `d1 >> 1;
		12'd356: toneL = `g1 >> 2;
		12'd357: toneL = `g1 >> 2;
		12'd358: toneL = `d1 >> 1;
		12'd359: toneL = `d1 >> 1;
		12'd360: toneL = `g1 >> 2;
		12'd361: toneL = `g1 >> 2;
		12'd362: toneL = `d1 >> 1;
		12'd363: toneL = `d1 >> 1;
		12'd364: toneL = `g1 >> 2;
		12'd365: toneL = `g1 >> 2;
		12'd366: toneL = `d1 >> 1;
		12'd367: toneL = `d1 >> 1;
		12'd368: toneL = `g1 >> 2;
		12'd369: toneL = `g1 >> 2;
		12'd370: toneL = `d1 >> 1;
		12'd371: toneL = `d1 >> 1;
		12'd372: toneL = `g1 >> 2;
		12'd373: toneL = `g1 >> 2;
		12'd374: toneL = `d1 >> 1;
		12'd375: toneL = `d1 >> 1;
		12'd376: toneL = `g1 >> 2;
		12'd377: toneL = `g1 >> 2;
		12'd378: toneL = `d1 >> 1;
		12'd379: toneL = `d1 >> 1;
		12'd380: toneL = `g1 >> 2;
		12'd381: toneL = `g1 >> 2;
		12'd382: toneL = `a1_d >> 2;
		12'd383: toneL = `a1_d >> 2;
		12'd384: toneL = `a1 >> 2;
		12'd385: toneL = `a1 >> 2;
		12'd386: toneL = `e1 >> 1;
		12'd387: toneL = `e1 >> 1;
		12'd388: toneL = `a1 >> 2;
		12'd389: toneL = `a1 >> 2;
		12'd390: toneL = `e1 >> 1;
		12'd391: toneL = `e1 >> 1;
		12'd392: toneL = `a1 >> 2;
		12'd393: toneL = `a1 >> 2;
		12'd394: toneL = `e1 >> 1;
		12'd395: toneL = `e1 >> 1;
		12'd396: toneL = `a1 >> 2;
		12'd397: toneL = `a1 >> 2;
		12'd398: toneL = `e1 >> 1;
		12'd399: toneL = `e1 >> 1;
		12'd400: toneL = `a1 >> 2;
		12'd401: toneL = `a1 >> 2;
		12'd402: toneL = `e1 >> 1;
		12'd403: toneL = `e1 >> 1;
		12'd404: toneL = `a1 >> 2;
		12'd405: toneL = `a1 >> 2;
		12'd406: toneL = `e1 >> 1;
		12'd407: toneL = `e1 >> 1;
		12'd408: toneL = `a1 >> 2;
		12'd409: toneL = `a1 >> 2;
		12'd410: toneL = `e1 >> 1;
		12'd411: toneL = `e1 >> 1;
		12'd412: toneL = `d1 >> 1;
		12'd413: toneL = `d1 >> 1;
		12'd414: toneL = `c1_u >> 1;
		12'd415: toneL = `c1_u >> 1;
		12'd416: toneL = `b1 >> 2;
		12'd417: toneL = `b1 >> 2;
		12'd418: toneL = `f1_u >> 1;
		12'd419: toneL = `f1_u >> 1;
		12'd420: toneL = `b1 >> 2;
		12'd421: toneL = `b1 >> 2;
		12'd422: toneL = `f1_u >> 1;
		12'd423: toneL = `f1_u >> 1;
		12'd424: toneL = `b1 >> 2;
		12'd425: toneL = `b1 >> 2;
		12'd426: toneL = `f1_u >> 1;
		12'd427: toneL = `f1_u >> 1;
		12'd428: toneL = `b1 >> 2;
		12'd429: toneL = `b1 >> 2;
		12'd430: toneL = `f1_u >> 1;
		12'd431: toneL = `f1_u >> 1;
		12'd432: toneL = `b1 >> 2;
		12'd433: toneL = `b1 >> 2;
		12'd434: toneL = `f1_u >> 1;
		12'd435: toneL = `f1_u >> 1;
		12'd436: toneL = `d1 >> 1;
		12'd437: toneL = `d1 >> 1;
		12'd438: toneL = `e1 >> 1;
		12'd439: toneL = `e1 >> 1;
		12'd440: toneL = `f1_u >> 1;
		12'd441: toneL = `f1_u >> 1;
		12'd442: toneL = `e1 >> 1;
		12'd443: toneL = `e1 >> 1;
		12'd444: toneL = `d1 >> 1;
		12'd445: toneL = `d1 >> 1;
		12'd446: toneL = `f1_u >> 1;
		12'd447: toneL = `f1_u >> 1;
		12'd448: toneL = `c1 >> 1;
		12'd449: toneL = `c1 >> 1;
		12'd450: toneL = `g1 >> 1;
		12'd451: toneL = `g1 >> 1;
		12'd452: toneL = `c1 >> 1;
		12'd453: toneL = `c1 >> 1;
		12'd454: toneL = `g1 >> 1;
		12'd455: toneL = `g1 >> 1;
		12'd456: toneL = `c1 >> 1;
		12'd457: toneL = `c1 >> 1;
		12'd458: toneL = `g1 >> 1;
		12'd459: toneL = `g1 >> 1;
		12'd460: toneL = `c1 >> 1;
		12'd461: toneL = `c1 >> 1;
		12'd462: toneL = `g1 >> 1;
		12'd463: toneL = `g1 >> 1;
		12'd464: toneL = `c1 >> 1;
		12'd465: toneL = `c1 >> 1;
		12'd466: toneL = `g1 >> 1;
		12'd467: toneL = `g1 >> 1;
		12'd468: toneL = `d1_u >> 1;
		12'd469: toneL = `d1_u >> 1;
		12'd470: toneL = `f1 >> 1;
		12'd471: toneL = `f1 >> 1;
		12'd472: toneL = `g1_d >> 1;
		12'd473: toneL = `g1_d >> 1;
		12'd474: toneL = `f1 >> 1;
		12'd475: toneL = `f1 >> 1;
		12'd476: toneL = `e1 >> 1;
		12'd477: toneL = `e1 >> 1;
		12'd478: toneL = `g1 >> 1;
		12'd479: toneL = `g1 >> 1;
		12'd480: toneL = `c1_u >> 1;
		12'd481: toneL = `c1_u >> 1;
		12'd482: toneL = `g1_u >> 1;
		12'd483: toneL = `g1_u >> 1;
		12'd484: toneL = `c1_u >> 1;
		12'd485: toneL = `c1_u >> 1;
		12'd486: toneL = `g1_u >> 1;
		12'd487: toneL = `g1_u >> 1;
		12'd488: toneL = `c1_u >> 1;
		12'd489: toneL = `c1_u >> 1;
		12'd490: toneL = `g1_u >> 1;
		12'd491: toneL = `g1_u >> 1;
		12'd492: toneL = `c1_u >> 1;
		12'd493: toneL = `c1_u >> 1;
		12'd494: toneL = `g1_u >> 1;
		12'd495: toneL = `g1_u >> 1;
		12'd496: toneL = `c1_u >> 1;
		12'd497: toneL = `c1_u >> 1;
		12'd498: toneL = `g1_u >> 1;
		12'd499: toneL = `g1_u >> 1;
		12'd500: toneL = `e1 >> 1;
		12'd501: toneL = `e1 >> 1;
		12'd502: toneL = `f1_u >> 1;
		12'd503: toneL = `f1_u >> 1;
		12'd504: toneL = `g1_u >> 1;
		12'd505: toneL = `g1_u >> 1;
		12'd506: toneL = `g1_d >> 1;
		12'd507: toneL = `g1_d >> 1;
		12'd508: toneL = `e1 >> 1;
		12'd509: toneL = `e1 >> 1;
		12'd510: toneL = `a1_d >> 1;
		12'd511: toneL = `a1_d >> 1;
		12'd512: toneL = `d1 >> 1;
		12'd513: toneL = `d1 >> 1;
		12'd514: toneL = `a1 >> 1;
		12'd515: toneL = `a1 >> 1;
		12'd516: toneL = `d1 >> 1;
		12'd517: toneL = `d1 >> 1;
		12'd518: toneL = `a1 >> 1;
		12'd519: toneL = `a1 >> 1;
		12'd520: toneL = `d1 >> 1;
		12'd521: toneL = `d1 >> 1;
		12'd522: toneL = `a1 >> 1;
		12'd523: toneL = `a1 >> 1;
		12'd524: toneL = `d1 >> 1;
		12'd525: toneL = `d1 >> 1;
		12'd526: toneL = `a1 >> 1;
		12'd527: toneL = `a1 >> 1;
		12'd528: toneL = `d1 >> 1;
		12'd529: toneL = `d1 >> 1;
		12'd530: toneL = `a1 >> 1;
		12'd531: toneL = `a1 >> 1;
		12'd532: toneL = `f1 >> 1;
		12'd533: toneL = `f1 >> 1;
		12'd534: toneL = `g1 >> 1;
		12'd535: toneL = `g1 >> 1;
		12'd536: toneL = `a1 >> 1;
		12'd537: toneL = `a1 >> 1;
		12'd538: toneL = `g1 >> 1;
		12'd539: toneL = `g1 >> 1;
		12'd540: toneL = `f1 >> 1;
		12'd541: toneL = `f1 >> 1;
		12'd542: toneL = `e1 >> 1;
		12'd543: toneL = `e1 >> 1;
		12'd544: toneL = `d1 >> 1;
		12'd545: toneL = `d1 >> 1;
		12'd546: toneL = `d1 >> 1;
		12'd547: toneL = `d1 >> 1;
		12'd548: toneL = `a1 >> 2;
		12'd549: toneL = `a1 >> 2;
		12'd550: toneL = `a1 >> 2;
		12'd551: toneL = `a1 >> 2;
		12'd552: toneL = `b1 >> 2;
		12'd553: toneL = `b1 >> 2;
		12'd554: toneL = `g1 >> 1;
		12'd555: toneL = `g1 >> 1;
		12'd556: toneL = `b1 >> 2;
		12'd557: toneL = `b1 >> 2;
		12'd558: toneL = `g1 >> 1;
		12'd559: toneL = `g1 >> 1;
		12'd560: toneL = `b1 >> 2;
		12'd561: toneL = `b1 >> 2;
		12'd562: toneL = `g1 >> 1;
		12'd563: toneL = `g1 >> 1;
		12'd564: toneL = `b1 >> 2;
		12'd565: toneL = `b1 >> 2;
		12'd566: toneL = `g1 >> 1;
		12'd567: toneL = `g1 >> 1;
		12'd568: toneL = `b1 >> 2;
		12'd569: toneL = `b1 >> 2;
		12'd570: toneL = `g1 >> 1;
		12'd571: toneL = `g1 >> 1;
		12'd572: toneL = `b1 >> 2;
		12'd573: toneL = `b1 >> 2;
		12'd574: toneL = `g1 >> 1;
		12'd575: toneL = `g1 >> 1;
		12'd576: toneL = `b1 >> 2;
		12'd577: toneL = `b1 >> 2;
		12'd578: toneL = `g1 >> 1;
		12'd579: toneL = `g1 >> 1;
		12'd580: toneL = `b1 >> 2;
		12'd581: toneL = `b1 >> 2;
		12'd582: toneL = `g1 >> 1;
		12'd583: toneL = `g1 >> 1;
		12'd584: toneL = `d1 >> 1;
		12'd585: toneL = `d1 >> 1;
		12'd586: toneL = `d1 >> 1;
		12'd587: toneL = `d1 >> 1;
		12'd588: toneL = `a1 >> 2;
		12'd589: toneL = `a1 >> 2;
		12'd590: toneL = `a1 >> 2;
		12'd591: toneL = `a1 >> 2;
		12'd592: toneL = `b1_d >> 2;
		12'd593: toneL = `b1_d >> 2;
		12'd594: toneL = `f1 >> 1;
		12'd595: toneL = `f1 >> 1;
		12'd596: toneL = `b1_d >> 2;
		12'd597: toneL = `b1_d >> 2;
		12'd598: toneL = `f1 >> 1;
		12'd599: toneL = `f1 >> 1;
		12'd600: toneL = `b1_d >> 2;
		12'd601: toneL = `b1_d >> 2;
		12'd602: toneL = `f1 >> 1;
		12'd603: toneL = `f1 >> 1;
		12'd604: toneL = `b1_d >> 2;
		12'd605: toneL = `b1_d >> 2;
		12'd606: toneL = `f1 >> 1;
		12'd607: toneL = `f1 >> 1;
		12'd608: toneL = `b1_d >> 2;
		12'd609: toneL = `b1_d >> 2;
		12'd610: toneL = `f1 >> 1;
		12'd611: toneL = `f1 >> 1;
		12'd612: toneL = `b1_d >> 2;
		12'd613: toneL = `b1_d >> 2;
		12'd614: toneL = `f1 >> 1;
		12'd615: toneL = `f1 >> 1;
		12'd616: toneL = `b1_d >> 2;
		12'd617: toneL = `b1_d >> 2;
		12'd618: toneL = `f1 >> 1;
		12'd619: toneL = `f1 >> 1;
		12'd620: toneL = `b1_d >> 2;
		12'd621: toneL = `b1_d >> 2;
		12'd622: toneL = `f1 >> 1;
		12'd623: toneL = `f1 >> 1;
		12'd624: toneL = `b1 >> 2;
		12'd625: toneL = `b1 >> 2;
		12'd626: toneL = `e1 >> 1;
		12'd627: toneL = `e1 >> 1;
		12'd628: toneL = `b1 >> 2;
		12'd629: toneL = `b1 >> 2;
		12'd630: toneL = `e1 >> 1;
		12'd631: toneL = `e1 >> 1;
		12'd632: toneL = `b1 >> 2;
		12'd633: toneL = `b1 >> 2;
		12'd634: toneL = `e1 >> 1;
		12'd635: toneL = `e1 >> 1;
		12'd636: toneL = `b1 >> 2;
		12'd637: toneL = `b1 >> 2;
		12'd638: toneL = `e1 >> 1;
		12'd639: toneL = `e1 >> 1;
		12'd640: toneL = `b1 >> 2;
		12'd641: toneL = `b1 >> 2;
		12'd642: toneL = `e1 >> 1;
		12'd643: toneL = `e1 >> 1;
		12'd644: toneL = `b1 >> 2;
		12'd645: toneL = `b1 >> 2;
		12'd646: toneL = `e1 >> 1;
		12'd647: toneL = `e1 >> 1;
		12'd648: toneL = `b1 >> 2;
		12'd649: toneL = `b1 >> 2;
		12'd650: toneL = `e1 >> 1;
		12'd651: toneL = `e1 >> 1;
		12'd652: toneL = `b1 >> 2;
		12'd653: toneL = `b1 >> 2;
		12'd654: toneL = `e1 >> 1;
		12'd655: toneL = `e1 >> 1;

		default : toneL = `non;
	endcase
end

always @ (*) begin
	if(pitch == 0) tone = toneH;
	else if(pitch == 1) tone = toneM;
	else if(pitch == 2) tone = toneL;
	else tone = toneM;
end


endmodule